 module forwarding_unit
	(
	);
	
	always@() begin
	end
endmodule
