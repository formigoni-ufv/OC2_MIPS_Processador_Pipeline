 module hazard_detection_unit
	(
	);
	
	always@() begin
	end
endmodule
